`include "types.sv"
